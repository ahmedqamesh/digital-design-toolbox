library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.std_logic_arith.all;
-- ===========================================================================
--  File: lab54.vhd
--  Author: Ahmed Qamesh
--  Date: 28/12/2025
-- ===========================================================================
--  Description: Pseudo random sequence generator from WiMAX and testbench for it. Perform simulations.
--  The delay block has two inputs (clocking and 8-bit width data) and one output (8-bit data word). 
-- ===========================================================================

entity lab54 is
    Port ( clk : in STD_LOGIC;
           srst : in STD_LOGIC;
           psp_bit : out STD_LOGIC);
end lab54;
architecture Behavioral of lab54 is

-- WiMAX stands for Worldwide Interoperability for Microwave Access
-- the standard defines pseudo-random sequences for scrambling and spreading signals.
-- These sequences are generated by linear feedback shift registers (LFSRs) based pseudo-random number generator (PRNG) 
-- The XOR of MSBs in the LFSR is directly part of WiMAX scrambling logic to randomize transmitted data.
signal lfsr : std_logic_vector(14 downto 0); -- 15-bit LFSR representing the WiMAX PRSG state.
signal xor_bit : std_logic; -- XOR of the two most significant bits
begin
-- XOR of MSB (bit 14) and next MSB (bit 13) calculated every cycle 
 xor_bit <= lfsr(14) xor lfsr(13);
process (clk) begin
	if rising_edge(clk) then
        if srst='1' then
        -- Initialize to 101010001110110
         lfsr <= "101010001110110";
        else
        -- Shift right with XOR feedback into LSB
        lfsr <= xor_bit & lfsr(14 downto 1);
        end if;
	end if;
end process;
 -- Output: XOR result immediately available
 psp_bit <= xor_bit;
end Behavioral;

